----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:25:04 10/04/2018 
-- Design Name: 
-- Module Name:    Decoder2_3 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Decoder2_3 is
    Port ( Sel : in  STD_LOGIC_VECTOR (1 DOWNTO 0);
           DEC : OUT STD_LOGIC_VECTOR (2 downto 0));
end Decoder2_3;

architecture Behavioral of Decoder2_3 is

begin

process (Sel)
begin
    DEC <= "111";        -- default output value
        case Sel is
            when "00" => DEC(0) <= '0';
            when "01" => DEC(1) <= '0';
            when "10" => DEC(2) <= '0';
            when others => DEC <= "111";
        end case;
end process;


end Behavioral;

